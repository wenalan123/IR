module  smg_decoder(
        input         [ 3: 0]  hex_in                   ,
        output  reg   [ 6: 0]  hex_out 
);
//=====================================================================\
// ********** Define Parameter and Internal Signals *************
//=====================================================================/



//======================================================================
// ***************      Main    Code    ****************
//======================================================================
//hex_out
always  @(*) begin
            case(hex_in)  //共阳极7段数码管，为低电平亮
                4'h0: hex_out     <=      7'b100_0000;                  
                4'h1: hex_out     <=      7'b111_1001;
                4'h2: hex_out     <=      7'b010_0100;
                4'h3: hex_out     <=      7'b011_0000;
                4'h4: hex_out     <=      7'b001_1001;
                4'h5: hex_out     <=      7'b001_0010;
                4'h6: hex_out     <=      7'b000_0010;
                4'h7: hex_out     <=      7'b111_1000;
                4'h8: hex_out     <=      7'b000_0000;
                4'h9: hex_out     <=      7'b001_0000;
                4'ha: hex_out     <=      7'b000_1000;
                4'hb: hex_out     <=      7'b000_0011;
                4'hc: hex_out     <=      7'b100_0110;
                4'hd: hex_out     <=      7'b010_0001;
                4'he: hex_out     <=      7'b000_0110;
                4'hf: hex_out     <=      7'b000_1110;

                default:
                      hex_out     <=      7'b100_0000;
            endcase
end



endmodule
